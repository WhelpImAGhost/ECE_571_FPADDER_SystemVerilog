//Module to Add Normalized Values Together

module ALU(fpbus.alu bus);



endmodule