module fpadder(fpbus);
 


endmodule